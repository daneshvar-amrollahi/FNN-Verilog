module bh_mem(
    bh0, bh1, bh2, bh3, bh4, bh5, bh6, bh7, bh8, bh9, bh10, bh11, bh12, bh13, bh14, bh15, 
    bh16, bh17, bh18, bh19, bh20, bh21, bh22, bh23, bh24, bh25, bh26, bh27, bh28, bh29;
);

    output [7 : 0] bh0, bh1, bh2, bh3, bh4, bh5, bh6, bh7, bh8, bh9, bh10, bh11, bh12, bh13, bh14, bh15, 
    bh16, bh17, bh18, bh19, bh20, bh21, bh22, bh23, bh24, bh25, bh26, bh27, bh28, bh29;


    assign bh0 = 8'b00110100;
    assign bh1 = 8'b00110110;
    assign bh2 = 8'b10010001;
    assign bh3 = 8'b11001110;
    assign bh4 = 8'b11110100;
    assign bh5 = 8'b11000111;
    assign bh6 = 8'b10011110;
    assign bh7 = 8'b11111111;
    assign bh8 = 8'b10111000;
    assign bh9 = 8'b11001111;
    assign bh10 = 8'b01000011;
    assign bh11 = 8'b11001001;
    assign bh12 = 8'b00010000;
    assign bh13 = 8'b00111001;
    assign bh14 = 8'b10110010;
    assign bh15 = 8'b11101010;
    assign bh16 = 8'b11010111;
    assign bh17 = 8'b11111111;
    assign bh18 = 8'b10011101;
    assign bh19 = 8'b10100001;
    assign bh20 = 8'b11101111;
    assign bh21 = 8'b01010011;
    assign bh22 = 8'b00100101;
    assign bh23 = 8'b11011100;
    assign bh24 = 8'b00101101;
    assign bh25 = 8'b10110110;
    assign bh26 = 8'b00001011;
    assign bh27 = 8'b11111011;
    assign bh28 = 8'b11111111;
    assign bh29 = 8'b11111111;

endmodule

endmodule