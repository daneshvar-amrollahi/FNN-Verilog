module wo_mem(
    wo0, wo1, wo2, wo3, wo4, wo5, wo6, wo7, wo8, wo9
);
    output [239 : 0] wo0, wo1, wo2, wo3, wo4, wo5, wo6, wo7, wo8, wo9;

    assign wo0 = 240'b00001100_10111010_10001010_10001101_10001010_10010000_10010000_00010001_00000001_00101111_00011101_00001100_00011001_10001011_00011101_10100011_10010111_10011110_10000001_00001011_00000011_10100100_10100111_10001110_00010101_00010000_00001101_10010101_00110110_10011001;
    assign wo1 = 240'b00110110_10100000_10000110_10001000_00000101_10001101_00000100_10000100_00011100_10100111_00010001_00100110_00001100_10101010_00011100_10001001_00111111_10100110_10101100_10010010_10000101_00000110_00101000_00001111_10011110_00011100_00001000_00001100_00011010_10000100;
    assign wo2 = 240'b10001101_10101000_10011111_00010111_10100101_00101000_10011010_00011111_10011110_00100010_00100100_00011101_00000110_00110101_10010001_10100110_10001110_00001011_10101101_10110110_00000100_10000011_10000111_10100101_10110010_10011000_10100010_00011110_10010010_10011110;
    assign wo3 = 240'b10111000_11011000_00000101_10001001_11001011_00001101_10101001_11001100_00000110_10100100_10101000_00001101_00000001_10101010_00011000_00111000_10100101_00100010_00000011_11001011_00011100_00000110_10000011_10000101_00010010_00001011_00000101_00011000_10000001_00001011;
    assign wo4 = 240'b10001101_00000011_10011001_00010001_00000100_10011010_10111011_10010000_10010001_01011010_10100011_11001100_01111010_10101110_00001101_10000101_00000011_10101101_10011011_00010001_10001101_10010011_00001001_10010100_10011100_10000110_10000111_00000100_10001000_10000010;
    assign wo5 = 240'b10111100_10010100_00000011_00100110_00110010_10100110_01010101_11100110_10000010_10101001_10010001_10011001_10101001_10000100_00001101_10111010_00010010_00001001_00110100_10011001_10010111_00111110_10000001_10011110_10111001_00101011_10011001_10000011_00001011_10000110;
    assign wo6 = 240'b00100001_10001000_00000110_10010111_00000001_00000001_00010101_00001010_00010000_10011101_10000100_00001110_10110100_00000111_10001011_10010001_10000011_00001111_00110110_00100110_00001011_00100011_00001101_00001100_00110000_00001110_00010111_10010101_10110001_10010011;
    assign wo7 = 240'b00010010_01110100_00101110_01010101_00100000_00001000_10000100_00101011_10011111_00000110_10101110_10011101_10110010_00000110_00001000_00010001_00001011_00001100_10000110_00010110_00000001_10010011_00010000_00011000_01000000_00010101_00000011_10011001_10000001_00000000;
    assign wo8 = 240'b10010101_11111111_10000011_10101010_00111111_10000010_10011011_00000010_10101010_00011011_10111011_10010111_10001011_00000001_10111110_10110001_10110110_10100001_10100000_00000001_10001000_10110000_10011001_00100110_10100011_10110110_10010010_10011111_10100011_00011110;
    assign wo9 = 240'b10101101_01111111_11101110_10101011_10101111_00001110_10011101_10111000_00010010_11111111_00001000_00001100_11110000_11010000_00001000_10000001_10011010_10010100_00010101_00001101_00000011_00100010_00010111_00001100_11011111_10001001_00001100_00001011_10001011_00000011;

endmodule